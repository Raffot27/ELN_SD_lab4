versione prova
